library ieee;
use ieee.std_logic_1164.all;

entity name is
port( variable1, varialbe2 : in std_logic;
		             variable3 : out std_logic);
end name;

architecture arc of name is
begin 

	q <= //boolean expressions;
	
end arc; 
